-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 10.1 Build 153 11/29/2010 SJ Full Version"
-- CREATED		"Fri Nov 18 19:06:39 2011"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Lab4_and_5 IS 
	PORT
	(
		InputA :  IN  STD_LOGIC;
		InputB :  IN  STD_LOGIC;
		InputC :  IN  STD_LOGIC;
		InputD :  IN  STD_LOGIC;
		OutputA :  OUT  STD_LOGIC;
		OutputB :  OUT  STD_LOGIC;
		OutputC :  OUT  STD_LOGIC;
		OutputD :  OUT  STD_LOGIC;
		OutputE :  OUT  STD_LOGIC;
		OutputF :  OUT  STD_LOGIC;
		OutputG :  OUT  STD_LOGIC
	);
END Lab4_and_5;

ARCHITECTURE bdf_type OF Lab4_and_5 IS 

SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_44 <= SYNTHESIZED_WIRE_65 AND InputB AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_50 <= SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND InputC AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_65 AND InputB AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_57 <= SYNTHESIZED_WIRE_65 AND InputB AND SYNTHESIZED_WIRE_67;


SYNTHESIZED_WIRE_58 <= InputA AND InputB AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_64 <= SYNTHESIZED_WIRE_65 AND InputB AND InputC AND InputD;


SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_65 AND InputB AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_47 <= InputB AND InputC AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_48 <= InputA AND InputB AND InputC;


SYNTHESIZED_WIRE_54 <= InputA AND SYNTHESIZED_WIRE_66 AND InputC AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_61 <= SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND InputD;


SYNTHESIZED_WIRE_62 <= InputA AND InputB AND SYNTHESIZED_WIRE_67 AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_41 <= InputA AND InputB AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_45 <= InputA AND InputB AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_49 <= InputA AND InputB AND SYNTHESIZED_WIRE_68;


SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67 AND InputD;


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_65 AND InputD;


SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND InputC;


SYNTHESIZED_WIRE_63 <= SYNTHESIZED_WIRE_65 AND SYNTHESIZED_WIRE_66 AND SYNTHESIZED_WIRE_67;


SYNTHESIZED_WIRE_42 <= InputA AND SYNTHESIZED_WIRE_66 AND InputC AND InputD;


SYNTHESIZED_WIRE_46 <= InputA AND InputC AND InputD;


SYNTHESIZED_WIRE_53 <= InputB AND InputC AND InputD;


SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_65 AND InputC AND InputD;


SYNTHESIZED_WIRE_65 <= NOT(InputA);



SYNTHESIZED_WIRE_66 <= NOT(InputB);



SYNTHESIZED_WIRE_67 <= NOT(InputC);



SYNTHESIZED_WIRE_68 <= NOT(InputD);



OutputA <= SYNTHESIZED_WIRE_40 OR SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42 OR SYNTHESIZED_WIRE_43;


OutputB <= SYNTHESIZED_WIRE_44 OR SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_46 OR SYNTHESIZED_WIRE_47;


OutputC <= SYNTHESIZED_WIRE_48 OR SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50;


OutputD <= SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_52 OR SYNTHESIZED_WIRE_53 OR SYNTHESIZED_WIRE_54;


OutputE <= SYNTHESIZED_WIRE_55 OR SYNTHESIZED_WIRE_56 OR SYNTHESIZED_WIRE_57;


OutputF <= SYNTHESIZED_WIRE_58 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_61;


OutputG <= SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_64;


END bdf_type;