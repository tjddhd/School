-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 10.1 Build 153 11/29/2010 SJ Full Version"
-- CREATED		"Wed Nov 16 14:18:27 2011"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Counter IS 
	PORT
	(
		InputX :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		RST :  IN  STD_LOGIC;
		OUTPUT1 :  OUT  STD_LOGIC;
		OUTPUT2 :  OUT  STD_LOGIC;
		OUTPUT3 :  OUT  STD_LOGIC
	);
END Counter;

ARCHITECTURE bdf_type OF Counter IS 

SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;


BEGIN 
OUTPUT1 <= SYNTHESIZED_WIRE_41;
OUTPUT2 <= SYNTHESIZED_WIRE_43;
OUTPUT3 <= SYNTHESIZED_WIRE_44;
SYNTHESIZED_WIRE_45 <= '1';



SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_35 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_41 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_41 AND InputX;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND InputX;


SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_41 AND InputX;


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43 AND InputX;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_44 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_41 AND InputX;


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_41;


SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_44 AND SYNTHESIZED_WIRE_38;


SYNTHESIZED_WIRE_36 <= SYNTHESIZED_WIRE_44 AND SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_40;


PROCESS(clk,RST,SYNTHESIZED_WIRE_45)
BEGIN
IF (RST = '0') THEN
	SYNTHESIZED_WIRE_44 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_44 <= SYNTHESIZED_WIRE_20;
END IF;
END PROCESS;


PROCESS(clk,RST,SYNTHESIZED_WIRE_45)
BEGIN
IF (RST = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_22;
END IF;
END PROCESS;


PROCESS(clk,RST,SYNTHESIZED_WIRE_45)
BEGIN
IF (RST = '0') THEN
	SYNTHESIZED_WIRE_41 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_41 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_24;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_39 <= NOT(SYNTHESIZED_WIRE_41);



SYNTHESIZED_WIRE_38 <= NOT(SYNTHESIZED_WIRE_43);



SYNTHESIZED_WIRE_42 <= NOT(SYNTHESIZED_WIRE_44);



SYNTHESIZED_WIRE_40 <= NOT(InputX);



SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27 OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_34 OR SYNTHESIZED_WIRE_35 OR SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37;


END bdf_type;